module top_module ( input a, input b, output out );
    mod_a top_module (a,b,out);
endmodule
