
// to write code for top module 

module top_module ( 
    input a, 
    input b, 
    input c,
    input d,
    output out1,
    output out2
);
   mod_a top_module (out1 , out2 , a, b, c, d);
endmodule
